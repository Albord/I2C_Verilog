/*
	Autor: Albert Espi�a Rojas
	Modulo: I2C_SLAVE_MEMORY
	Modulo de memoria. Podemos acceder y guardar datos. 
	El modulo tiene como parametro, el tama�o de la direcci�n de memoria, el n�mero de direcci�nes ,es decir el n�mero de datos
	y el n�mero de bytes en los datos

*/

module I2C_SLAVE_MEMORY #( parameter ADDRESSLENGTH, parameter ADDRESSNUM, parameter NBYTES)(Enable, RorW, DirectionBuffer, InputBuffer, OutputBuffer, AddressFound, AddressList);
	input Enable; //
	input RorW;
	input [((ADDRESSLENGTH)*ADDRESSNUM) - 1: 0]AddressList;
	output reg AddressFound = 1'b0;
	input wire [(ADDRESSLENGTH-1): 0] DirectionBuffer;
	input wire [7:0]InputBuffer;
	output reg [7:0]OutputBuffer;
	reg [8*NBYTES*ADDRESSNUM: 0 ] Data = 1'b0;
	integer LocalAddressID = 0;
	integer ByteCounter = 0;
	

always @(posedge Enable)//Si se activa el enable, es cuando transferimos los datos del buffer a la memoria
begin
	 //Modo transferencia, intercambiamos datos entre el buffer y los datos de la memoria
	if (RorW) Data[LocalAddressID*8*NBYTES + (ByteCounter)*(8) +:8] <= InputBuffer;
	else OutputBuffer <= Data[LocalAddressID*8*NBYTES + (ByteCounter)*(8) +:8];
	if (ByteCounter < NBYTES - 1) ByteCounter <= ByteCounter + 1;
	else ByteCounter <= 0;
end

always@(DirectionBuffer) begin
	AddressFound = 1'b0;
	ByteCounter = 0;
	LocalAddressID = 0;
	for(LocalAddressID = 0; (LocalAddressID < ADDRESSNUM) &&  !AddressFound; LocalAddressID = LocalAddressID + 1) begin
		if (AddressList[ADDRESSLENGTH*(LocalAddressID)+:8] == DirectionBuffer) AddressFound = 1'b1;
	end
end


endmodule